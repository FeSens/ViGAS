// god_bless_apollo.v

// Generated using ACDS version 14.1 190 at 2015.06.02.11:06:06

`timescale 1 ps / 1 ps
module god_bless_apollo (
		input  wire        clk_clk,              //      clk.clk
		output wire [14:0] memory_mem_a,         //   memory.mem_a
		output wire [2:0]  memory_mem_ba,        //         .mem_ba
		output wire [0:0]  memory_mem_ck,        //         .mem_ck
		output wire [0:0]  memory_mem_ck_n,      //         .mem_ck_n
		output wire [0:0]  memory_mem_cke,       //         .mem_cke
		output wire [0:0]  memory_mem_cs_n,      //         .mem_cs_n
		output wire [3:0]  memory_mem_dm,        //         .mem_dm
		output wire [0:0]  memory_mem_ras_n,     //         .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,     //         .mem_cas_n
		output wire [0:0]  memory_mem_we_n,      //         .mem_we_n
		output wire        memory_mem_reset_n,   //         .mem_reset_n
		inout  wire [31:0] memory_mem_dq,        //         .mem_dq
		inout  wire [3:0]  memory_mem_dqs,       //         .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,     //         .mem_dqs_n
		output wire [0:0]  memory_mem_odt,       //         .mem_odt
		output wire [12:0] memory_0_mem_a,       // memory_0.mem_a
		output wire [2:0]  memory_0_mem_ba,      //         .mem_ba
		output wire        memory_0_mem_ck,      //         .mem_ck
		output wire        memory_0_mem_ck_n,    //         .mem_ck_n
		output wire        memory_0_mem_cke,     //         .mem_cke
		output wire        memory_0_mem_cs_n,    //         .mem_cs_n
		output wire        memory_0_mem_ras_n,   //         .mem_ras_n
		output wire        memory_0_mem_cas_n,   //         .mem_cas_n
		output wire        memory_0_mem_we_n,    //         .mem_we_n
		output wire        memory_0_mem_reset_n, //         .mem_reset_n
		inout  wire [7:0]  memory_0_mem_dq,      //         .mem_dq
		inout  wire        memory_0_mem_dqs,     //         .mem_dqs
		inout  wire        memory_0_mem_dqs_n,   //         .mem_dqs_n
		output wire        memory_0_mem_odt,     //         .mem_odt
		output wire        memory_0_mem_dm,      //         .mem_dm
		input  wire        memory_0_oct_rzqin,   //         .oct_rzqin
		input  wire        oct_rzqin,            //      oct.rzqin
		input  wire        reset_reset_n,        //    reset.reset_n
		output wire [7:0]  vga_red,              //      vga.red
		output wire [7:0]  vga_green,            //         .green
		output wire [7:0]  vga_blue,             //         .blue
		output wire        vga_hs,               //         .hs
		output wire        vga_vs,               //         .vs
		output wire        vga_sync,             //         .sync
		output wire        vga_blank,            //         .blank
		input  wire [3:0]  vga_sw,               //         .sw
		output wire        vga_clk_clk           //  vga_clk.clk
	);

	wire         pll_0_outclk0_clk;                                             // pll_0:outclk_0 -> Apollo_VIdeo_Processment_Unit_0:clk_25
	wire         pll_0_outclk1_clk;                                             // pll_0:outclk_1 -> [Apollo_VIdeo_Processment_Unit_0:clk_Avalon, hps_0:h2f_axi_clk, mem_if_ddr3_emif_0:mp_cmd_clk_0_clk, mem_if_ddr3_emif_0:mp_cmd_clk_1_clk, mem_if_ddr3_emif_0:mp_rfifo_clk_0_clk, mem_if_ddr3_emif_0:mp_rfifo_clk_1_clk, mem_if_ddr3_emif_0:mp_wfifo_clk_0_clk, mem_if_ddr3_emif_0:mp_wfifo_clk_1_clk, mm_interconnect_0:pll_0_outclk1_clk, mm_interconnect_1:pll_0_outclk1_clk, rst_controller_001:clk, rst_controller_002:clk]
	wire  [31:0] apollo_video_processment_unit_0_avalon_master_readdata;        // mm_interconnect_0:Apollo_VIdeo_Processment_Unit_0_avalon_master_readdata -> Apollo_VIdeo_Processment_Unit_0:read_readdata
	wire         apollo_video_processment_unit_0_avalon_master_waitrequest;     // mm_interconnect_0:Apollo_VIdeo_Processment_Unit_0_avalon_master_waitrequest -> Apollo_VIdeo_Processment_Unit_0:read_waitrequest
	wire         apollo_video_processment_unit_0_avalon_master_read;            // Apollo_VIdeo_Processment_Unit_0:read_request -> mm_interconnect_0:Apollo_VIdeo_Processment_Unit_0_avalon_master_read
	wire  [31:0] apollo_video_processment_unit_0_avalon_master_address;         // Apollo_VIdeo_Processment_Unit_0:read_address -> mm_interconnect_0:Apollo_VIdeo_Processment_Unit_0_avalon_master_address
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer; // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin_0
	wire  [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata;           // mem_if_ddr3_emif_0:avl_rdata_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_readdata
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest;        // mem_if_ddr3_emif_0:avl_ready_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_waitrequest
	wire  [27:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address;            // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_address -> mem_if_ddr3_emif_0:avl_addr_0
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read;               // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_read -> mem_if_ddr3_emif_0:avl_read_req_0
	wire   [3:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_byteenable -> mem_if_ddr3_emif_0:avl_be_0
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid;      // mem_if_ddr3_emif_0:avl_rdata_valid_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_readdatavalid
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write;              // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_write -> mem_if_ddr3_emif_0:avl_write_req_0
	wire  [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata;          // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_writedata -> mem_if_ddr3_emif_0:avl_wdata_0
	wire   [2:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_burstcount -> mem_if_ddr3_emif_0:avl_size_0
	wire   [1:0] hps_0_h2f_axi_master_awburst;                                  // hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                                    // hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                                    // hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                                   // mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                                      // mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                                   // hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                                    // hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                                      // hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                                  // hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                                   // hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                                   // hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                                   // hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                                   // hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	wire  [31:0] hps_0_h2f_axi_master_wdata;                                    // hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                                  // hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                                  // hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                                     // hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                                   // hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                                   // hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                                   // hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                                    // mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                                  // mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [31:0] hps_0_h2f_axi_master_rdata;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                                  // mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                                  // hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                                   // hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                                   // hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                                    // hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                                     // hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                                      // mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                                   // mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                                   // hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                                  // hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                                   // mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_beginbursttransfer; // mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin_1
	wire  [31:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_readdata;           // mem_if_ddr3_emif_0:avl_rdata_1 -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_readdata
	wire         mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_waitrequest;        // mem_if_ddr3_emif_0:avl_ready_1 -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_waitrequest
	wire  [27:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_address;            // mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_address -> mem_if_ddr3_emif_0:avl_addr_1
	wire         mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_read;               // mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_read -> mem_if_ddr3_emif_0:avl_read_req_1
	wire   [3:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_byteenable;         // mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_byteenable -> mem_if_ddr3_emif_0:avl_be_1
	wire         mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_readdatavalid;      // mem_if_ddr3_emif_0:avl_rdata_valid_1 -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_readdatavalid
	wire         mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_write;              // mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_write -> mem_if_ddr3_emif_0:avl_write_req_1
	wire  [31:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_writedata;          // mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_writedata -> mem_if_ddr3_emif_0:avl_wdata_1
	wire   [2:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_burstcount;         // mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_burstcount -> mem_if_ddr3_emif_0:avl_size_1
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> Apollo_VIdeo_Processment_Unit_0:reset
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [mm_interconnect_0:Apollo_VIdeo_Processment_Unit_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset, mm_interconnect_1:mem_if_ddr3_emif_0_avl_1_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mem_if_ddr3_emif_0_mp_cmd_reset_n_1_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                                         // hps_0:h2f_rst_n -> rst_controller_002:reset_in0

	Vga apollo_video_processment_unit_0 (
		.clk              (clk_clk),                                                   //         clock.clk
		.reset            (rst_controller_reset_out_reset),                            //         reset.reset
		.read_request     (apollo_video_processment_unit_0_avalon_master_read),        // avalon_master.read
		.read_address     (apollo_video_processment_unit_0_avalon_master_address),     //              .address
		.read_readdata    (apollo_video_processment_unit_0_avalon_master_readdata),    //              .readdata
		.read_waitrequest (apollo_video_processment_unit_0_avalon_master_waitrequest), //              .waitrequest
		.clk_25           (pll_0_outclk0_clk),                                         //        clk_25.clk
		.VGA_CLK          (vga_clk_clk),                                               //       VGA_clk.clk
		.VGA_R            (vga_red),                                                   //           VGA.red
		.VGA_G            (vga_green),                                                 //              .green
		.VGA_B            (vga_blue),                                                  //              .blue
		.VGA_HS           (vga_hs),                                                    //              .hs
		.VGA_VS           (vga_vs),                                                    //              .vs
		.VGA_SYNC_n       (vga_sync),                                                  //              .sync
		.VGA_BLANK_n      (vga_blank),                                                 //              .blank
		.sw               (vga_sw),                                                    //              .sw
		.clk_Avalon       (pll_0_outclk1_clk)                                          //  clock_Avalon.clk
	);

	god_bless_apollo_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a       (memory_0_mem_a),               //         memory.mem_a
		.mem_ba      (memory_0_mem_ba),              //               .mem_ba
		.mem_ck      (memory_0_mem_ck),              //               .mem_ck
		.mem_ck_n    (memory_0_mem_ck_n),            //               .mem_ck_n
		.mem_cke     (memory_0_mem_cke),             //               .mem_cke
		.mem_cs_n    (memory_0_mem_cs_n),            //               .mem_cs_n
		.mem_ras_n   (memory_0_mem_ras_n),           //               .mem_ras_n
		.mem_cas_n   (memory_0_mem_cas_n),           //               .mem_cas_n
		.mem_we_n    (memory_0_mem_we_n),            //               .mem_we_n
		.mem_reset_n (memory_0_mem_reset_n),         //               .mem_reset_n
		.mem_dq      (memory_0_mem_dq),              //               .mem_dq
		.mem_dqs     (memory_0_mem_dqs),             //               .mem_dqs
		.mem_dqs_n   (memory_0_mem_dqs_n),           //               .mem_dqs_n
		.mem_odt     (memory_0_mem_odt),             //               .mem_odt
		.mem_dm      (memory_0_mem_dm),              //               .mem_dm
		.oct_rzqin   (memory_0_oct_rzqin),           //               .oct_rzqin
		.h2f_rst_n   (hps_0_h2f_reset_reset),        //      h2f_reset.reset_n
		.h2f_axi_clk (pll_0_outclk1_clk),            //  h2f_axi_clock.clk
		.h2f_AWID    (hps_0_h2f_axi_master_awid),    // h2f_axi_master.awid
		.h2f_AWADDR  (hps_0_h2f_axi_master_awaddr),  //               .awaddr
		.h2f_AWLEN   (hps_0_h2f_axi_master_awlen),   //               .awlen
		.h2f_AWSIZE  (hps_0_h2f_axi_master_awsize),  //               .awsize
		.h2f_AWBURST (hps_0_h2f_axi_master_awburst), //               .awburst
		.h2f_AWLOCK  (hps_0_h2f_axi_master_awlock),  //               .awlock
		.h2f_AWCACHE (hps_0_h2f_axi_master_awcache), //               .awcache
		.h2f_AWPROT  (hps_0_h2f_axi_master_awprot),  //               .awprot
		.h2f_AWVALID (hps_0_h2f_axi_master_awvalid), //               .awvalid
		.h2f_AWREADY (hps_0_h2f_axi_master_awready), //               .awready
		.h2f_WID     (hps_0_h2f_axi_master_wid),     //               .wid
		.h2f_WDATA   (hps_0_h2f_axi_master_wdata),   //               .wdata
		.h2f_WSTRB   (hps_0_h2f_axi_master_wstrb),   //               .wstrb
		.h2f_WLAST   (hps_0_h2f_axi_master_wlast),   //               .wlast
		.h2f_WVALID  (hps_0_h2f_axi_master_wvalid),  //               .wvalid
		.h2f_WREADY  (hps_0_h2f_axi_master_wready),  //               .wready
		.h2f_BID     (hps_0_h2f_axi_master_bid),     //               .bid
		.h2f_BRESP   (hps_0_h2f_axi_master_bresp),   //               .bresp
		.h2f_BVALID  (hps_0_h2f_axi_master_bvalid),  //               .bvalid
		.h2f_BREADY  (hps_0_h2f_axi_master_bready),  //               .bready
		.h2f_ARID    (hps_0_h2f_axi_master_arid),    //               .arid
		.h2f_ARADDR  (hps_0_h2f_axi_master_araddr),  //               .araddr
		.h2f_ARLEN   (hps_0_h2f_axi_master_arlen),   //               .arlen
		.h2f_ARSIZE  (hps_0_h2f_axi_master_arsize),  //               .arsize
		.h2f_ARBURST (hps_0_h2f_axi_master_arburst), //               .arburst
		.h2f_ARLOCK  (hps_0_h2f_axi_master_arlock),  //               .arlock
		.h2f_ARCACHE (hps_0_h2f_axi_master_arcache), //               .arcache
		.h2f_ARPROT  (hps_0_h2f_axi_master_arprot),  //               .arprot
		.h2f_ARVALID (hps_0_h2f_axi_master_arvalid), //               .arvalid
		.h2f_ARREADY (hps_0_h2f_axi_master_arready), //               .arready
		.h2f_RID     (hps_0_h2f_axi_master_rid),     //               .rid
		.h2f_RDATA   (hps_0_h2f_axi_master_rdata),   //               .rdata
		.h2f_RRESP   (hps_0_h2f_axi_master_rresp),   //               .rresp
		.h2f_RLAST   (hps_0_h2f_axi_master_rlast),   //               .rlast
		.h2f_RVALID  (hps_0_h2f_axi_master_rvalid),  //               .rvalid
		.h2f_RREADY  (hps_0_h2f_axi_master_rready)   //               .rready
	);

	god_bless_apollo_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk                (clk_clk),                                                       //        pll_ref_clk.clk
		.global_reset_n             (reset_reset_n),                                                 //       global_reset.reset_n
		.soft_reset_n               (reset_reset_n),                                                 //         soft_reset.reset_n
		.afi_clk                    (),                                                              //            afi_clk.clk
		.afi_half_clk               (),                                                              //       afi_half_clk.clk
		.afi_reset_n                (),                                                              //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                              //   afi_reset_export.reset_n
		.mem_a                      (memory_mem_a),                                                  //             memory.mem_a
		.mem_ba                     (memory_mem_ba),                                                 //                   .mem_ba
		.mem_ck                     (memory_mem_ck),                                                 //                   .mem_ck
		.mem_ck_n                   (memory_mem_ck_n),                                               //                   .mem_ck_n
		.mem_cke                    (memory_mem_cke),                                                //                   .mem_cke
		.mem_cs_n                   (memory_mem_cs_n),                                               //                   .mem_cs_n
		.mem_dm                     (memory_mem_dm),                                                 //                   .mem_dm
		.mem_ras_n                  (memory_mem_ras_n),                                              //                   .mem_ras_n
		.mem_cas_n                  (memory_mem_cas_n),                                              //                   .mem_cas_n
		.mem_we_n                   (memory_mem_we_n),                                               //                   .mem_we_n
		.mem_reset_n                (memory_mem_reset_n),                                            //                   .mem_reset_n
		.mem_dq                     (memory_mem_dq),                                                 //                   .mem_dq
		.mem_dqs                    (memory_mem_dqs),                                                //                   .mem_dqs
		.mem_dqs_n                  (memory_mem_dqs_n),                                              //                   .mem_dqs_n
		.mem_odt                    (memory_mem_odt),                                                //                   .mem_odt
		.avl_ready_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest),        //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_0                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address),            //                   .address
		.avl_rdata_valid_0          (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid),      //                   .readdatavalid
		.avl_rdata_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata),           //                   .readdata
		.avl_wdata_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata),          //                   .writedata
		.avl_be_0                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable),         //                   .byteenable
		.avl_read_req_0             (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read),               //                   .read
		.avl_write_req_0            (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write),              //                   .write
		.avl_size_0                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount),         //                   .burstcount
		.avl_ready_1                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_waitrequest),        //              avl_1.waitrequest_n
		.avl_burstbegin_1           (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_1                 (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_address),            //                   .address
		.avl_rdata_valid_1          (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_readdatavalid),      //                   .readdatavalid
		.avl_rdata_1                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_readdata),           //                   .readdata
		.avl_wdata_1                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_writedata),          //                   .writedata
		.avl_be_1                   (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_byteenable),         //                   .byteenable
		.avl_read_req_1             (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_read),               //                   .read
		.avl_write_req_1            (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_write),              //                   .write
		.avl_size_1                 (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_burstcount),         //                   .burstcount
		.mp_cmd_clk_0_clk           (pll_0_outclk1_clk),                                             //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (reset_reset_n),                                                 //   mp_cmd_reset_n_0.reset_n
		.mp_cmd_clk_1_clk           (pll_0_outclk1_clk),                                             //       mp_cmd_clk_1.clk
		.mp_cmd_reset_n_1_reset_n   (reset_reset_n),                                                 //   mp_cmd_reset_n_1.reset_n
		.mp_rfifo_clk_0_clk         (pll_0_outclk1_clk),                                             //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (reset_reset_n),                                                 // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (pll_0_outclk1_clk),                                             //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (reset_reset_n),                                                 // mp_wfifo_reset_n_0.reset_n
		.mp_rfifo_clk_1_clk         (pll_0_outclk1_clk),                                             //     mp_rfifo_clk_1.clk
		.mp_rfifo_reset_n_1_reset_n (reset_reset_n),                                                 // mp_rfifo_reset_n_1.reset_n
		.mp_wfifo_clk_1_clk         (pll_0_outclk1_clk),                                             //     mp_wfifo_clk_1.clk
		.mp_wfifo_reset_n_1_reset_n (reset_reset_n),                                                 // mp_wfifo_reset_n_1.reset_n
		.local_init_done            (),                                                              //             status.local_init_done
		.local_cal_success          (),                                                              //                   .local_cal_success
		.local_cal_fail             (),                                                              //                   .local_cal_fail
		.oct_rzqin                  (oct_rzqin),                                                     //                oct.rzqin
		.pll_mem_clk                (),                                                              //        pll_sharing.pll_mem_clk
		.pll_write_clk              (),                                                              //                   .pll_write_clk
		.pll_locked                 (),                                                              //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (),                                                              //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (),                                                              //                   .pll_addr_cmd_clk
		.pll_avl_clk                (),                                                              //                   .pll_avl_clk
		.pll_config_clk             (),                                                              //                   .pll_config_clk
		.pll_mem_phy_clk            (),                                                              //                   .pll_mem_phy_clk
		.afi_phy_clk                (),                                                              //                   .afi_phy_clk
		.pll_avl_phy_clk            ()                                                               //                   .pll_avl_phy_clk
	);

	god_bless_apollo_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk), // outclk1.clk
		.locked   ()                   //  locked.export
	);

	god_bless_apollo_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk1_clk                                                 (pll_0_outclk1_clk),                                             //                                               pll_0_outclk1.clk
		.Apollo_VIdeo_Processment_Unit_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                            // Apollo_VIdeo_Processment_Unit_0_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),                            //   mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
		.Apollo_VIdeo_Processment_Unit_0_avalon_master_address             (apollo_video_processment_unit_0_avalon_master_address),         //               Apollo_VIdeo_Processment_Unit_0_avalon_master.address
		.Apollo_VIdeo_Processment_Unit_0_avalon_master_waitrequest         (apollo_video_processment_unit_0_avalon_master_waitrequest),     //                                                            .waitrequest
		.Apollo_VIdeo_Processment_Unit_0_avalon_master_read                (apollo_video_processment_unit_0_avalon_master_read),            //                                                            .read
		.Apollo_VIdeo_Processment_Unit_0_avalon_master_readdata            (apollo_video_processment_unit_0_avalon_master_readdata),        //                                                            .readdata
		.mem_if_ddr3_emif_0_avl_0_address                                  (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address),            //                                    mem_if_ddr3_emif_0_avl_0.address
		.mem_if_ddr3_emif_0_avl_0_write                                    (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write),              //                                                            .write
		.mem_if_ddr3_emif_0_avl_0_read                                     (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read),               //                                                            .read
		.mem_if_ddr3_emif_0_avl_0_readdata                                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata),           //                                                            .readdata
		.mem_if_ddr3_emif_0_avl_0_writedata                                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata),          //                                                            .writedata
		.mem_if_ddr3_emif_0_avl_0_beginbursttransfer                       (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer), //                                                            .beginbursttransfer
		.mem_if_ddr3_emif_0_avl_0_burstcount                               (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount),         //                                                            .burstcount
		.mem_if_ddr3_emif_0_avl_0_byteenable                               (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable),         //                                                            .byteenable
		.mem_if_ddr3_emif_0_avl_0_readdatavalid                            (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid),      //                                                            .readdatavalid
		.mem_if_ddr3_emif_0_avl_0_waitrequest                              (~mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest)        //                                                            .waitrequest
	);

	god_bless_apollo_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_axi_master_awid                                             (hps_0_h2f_axi_master_awid),                                     //                                            hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                           (hps_0_h2f_axi_master_awaddr),                                   //                                                                .awaddr
		.hps_0_h2f_axi_master_awlen                                            (hps_0_h2f_axi_master_awlen),                                    //                                                                .awlen
		.hps_0_h2f_axi_master_awsize                                           (hps_0_h2f_axi_master_awsize),                                   //                                                                .awsize
		.hps_0_h2f_axi_master_awburst                                          (hps_0_h2f_axi_master_awburst),                                  //                                                                .awburst
		.hps_0_h2f_axi_master_awlock                                           (hps_0_h2f_axi_master_awlock),                                   //                                                                .awlock
		.hps_0_h2f_axi_master_awcache                                          (hps_0_h2f_axi_master_awcache),                                  //                                                                .awcache
		.hps_0_h2f_axi_master_awprot                                           (hps_0_h2f_axi_master_awprot),                                   //                                                                .awprot
		.hps_0_h2f_axi_master_awvalid                                          (hps_0_h2f_axi_master_awvalid),                                  //                                                                .awvalid
		.hps_0_h2f_axi_master_awready                                          (hps_0_h2f_axi_master_awready),                                  //                                                                .awready
		.hps_0_h2f_axi_master_wid                                              (hps_0_h2f_axi_master_wid),                                      //                                                                .wid
		.hps_0_h2f_axi_master_wdata                                            (hps_0_h2f_axi_master_wdata),                                    //                                                                .wdata
		.hps_0_h2f_axi_master_wstrb                                            (hps_0_h2f_axi_master_wstrb),                                    //                                                                .wstrb
		.hps_0_h2f_axi_master_wlast                                            (hps_0_h2f_axi_master_wlast),                                    //                                                                .wlast
		.hps_0_h2f_axi_master_wvalid                                           (hps_0_h2f_axi_master_wvalid),                                   //                                                                .wvalid
		.hps_0_h2f_axi_master_wready                                           (hps_0_h2f_axi_master_wready),                                   //                                                                .wready
		.hps_0_h2f_axi_master_bid                                              (hps_0_h2f_axi_master_bid),                                      //                                                                .bid
		.hps_0_h2f_axi_master_bresp                                            (hps_0_h2f_axi_master_bresp),                                    //                                                                .bresp
		.hps_0_h2f_axi_master_bvalid                                           (hps_0_h2f_axi_master_bvalid),                                   //                                                                .bvalid
		.hps_0_h2f_axi_master_bready                                           (hps_0_h2f_axi_master_bready),                                   //                                                                .bready
		.hps_0_h2f_axi_master_arid                                             (hps_0_h2f_axi_master_arid),                                     //                                                                .arid
		.hps_0_h2f_axi_master_araddr                                           (hps_0_h2f_axi_master_araddr),                                   //                                                                .araddr
		.hps_0_h2f_axi_master_arlen                                            (hps_0_h2f_axi_master_arlen),                                    //                                                                .arlen
		.hps_0_h2f_axi_master_arsize                                           (hps_0_h2f_axi_master_arsize),                                   //                                                                .arsize
		.hps_0_h2f_axi_master_arburst                                          (hps_0_h2f_axi_master_arburst),                                  //                                                                .arburst
		.hps_0_h2f_axi_master_arlock                                           (hps_0_h2f_axi_master_arlock),                                   //                                                                .arlock
		.hps_0_h2f_axi_master_arcache                                          (hps_0_h2f_axi_master_arcache),                                  //                                                                .arcache
		.hps_0_h2f_axi_master_arprot                                           (hps_0_h2f_axi_master_arprot),                                   //                                                                .arprot
		.hps_0_h2f_axi_master_arvalid                                          (hps_0_h2f_axi_master_arvalid),                                  //                                                                .arvalid
		.hps_0_h2f_axi_master_arready                                          (hps_0_h2f_axi_master_arready),                                  //                                                                .arready
		.hps_0_h2f_axi_master_rid                                              (hps_0_h2f_axi_master_rid),                                      //                                                                .rid
		.hps_0_h2f_axi_master_rdata                                            (hps_0_h2f_axi_master_rdata),                                    //                                                                .rdata
		.hps_0_h2f_axi_master_rresp                                            (hps_0_h2f_axi_master_rresp),                                    //                                                                .rresp
		.hps_0_h2f_axi_master_rlast                                            (hps_0_h2f_axi_master_rlast),                                    //                                                                .rlast
		.hps_0_h2f_axi_master_rvalid                                           (hps_0_h2f_axi_master_rvalid),                                   //                                                                .rvalid
		.hps_0_h2f_axi_master_rready                                           (hps_0_h2f_axi_master_rready),                                   //                                                                .rready
		.pll_0_outclk1_clk                                                     (pll_0_outclk1_clk),                                             //                                                   pll_0_outclk1.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset      (rst_controller_002_reset_out_reset),                            //      hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_avl_1_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                            // mem_if_ddr3_emif_0_avl_1_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_mp_cmd_reset_n_1_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                            //       mem_if_ddr3_emif_0_mp_cmd_reset_n_1_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_avl_1_address                                      (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_address),            //                                        mem_if_ddr3_emif_0_avl_1.address
		.mem_if_ddr3_emif_0_avl_1_write                                        (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_write),              //                                                                .write
		.mem_if_ddr3_emif_0_avl_1_read                                         (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_read),               //                                                                .read
		.mem_if_ddr3_emif_0_avl_1_readdata                                     (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_readdata),           //                                                                .readdata
		.mem_if_ddr3_emif_0_avl_1_writedata                                    (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_writedata),          //                                                                .writedata
		.mem_if_ddr3_emif_0_avl_1_beginbursttransfer                           (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_beginbursttransfer), //                                                                .beginbursttransfer
		.mem_if_ddr3_emif_0_avl_1_burstcount                                   (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_burstcount),         //                                                                .burstcount
		.mem_if_ddr3_emif_0_avl_1_byteenable                                   (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_byteenable),         //                                                                .byteenable
		.mem_if_ddr3_emif_0_avl_1_readdatavalid                                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_readdatavalid),      //                                                                .readdatavalid
		.mem_if_ddr3_emif_0_avl_1_waitrequest                                  (~mm_interconnect_1_mem_if_ddr3_emif_0_avl_1_waitrequest)        //                                                                .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk1_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (pll_0_outclk1_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
